module unidadcontrol(input wire clk, reset, wez input wire [5:0] Opcode, output wire s_inc, s_inm_ we, wez, output wire [2:0] ;)

endmodule